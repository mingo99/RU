module ru #(
    parameter COL = 8
) (
    //verilog_format: off
    input clk,rstn
    //verilog_format: on
);

endmodule
